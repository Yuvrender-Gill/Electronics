module score();
endmodule 