module collision();
endmodule 