module enemy();
endmodule 