module healthKit();
endmodule 