module health();
endmodule 