module target();
endmodule 