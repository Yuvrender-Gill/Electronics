module enemyTop();
endmodule 