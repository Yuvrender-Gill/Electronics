module horribleEnemy();
endmodule 