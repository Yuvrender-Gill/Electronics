module gameLogo():
endmodule 