module gameFSM();
endmodule 