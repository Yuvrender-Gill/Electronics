module enemyBottom();
endmodule 