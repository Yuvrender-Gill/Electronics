module gameOver();
endmodule 