module grounded();
endmodule 