module keyboard_controller();
endmodule 